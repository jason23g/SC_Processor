-------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-------------------------------------------------------------------------------
ENTITY ALU_TB IS
END ALU_TB;
-------------------------------------------------------------------------------
ARCHITECTURE behavior OF ALU_TB IS

	-- Component Declaration for the Unit Under Test (UUT)

	COMPONENT ALU
	PORT (
		A		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		B		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Op		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Cout	: OUT STD_LOGIC;
		Zero	: OUT STD_LOGIC;
		Ovf		: OUT STD_LOGIC;
		Output	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
	END COMPONENT;

	--Inputs
	SIGNAL A	: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL B	: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Op	: STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
	
	--Outputs
	SIGNAL Cout		: STD_LOGIC;
	SIGNAL Zero		: STD_LOGIC;
	SIGNAL Ovf		: STD_LOGIC;
	SIGNAL Output	: STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	-- Instantiate the Unit Under Test (UUT)
	uut : ALU
	PORT MAP (
		A		=> A, 
		B		=> B, 
		Op		=> Op, 
		Cout	=> Cout, 
		Zero	=> Zero, 
		Ovf		=> Ovf, 
		Output	=> Output
	);
	
	-- Stimulus process
	stim_proc : PROCESS
	BEGIN
--		--------------- Addition --------------
--		Op <= "0000";--Add_1
--		A <= "00000000000000000000000000000000";
--		B <= "00000000000000000000000000000000";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_2
--		A <= "00000000001100001111100000011001";
--		B <= "00000001111100011001110000010001";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_3
--		A <= "00000000001100001111100000011001";
--		B <= "10000001111100011001110000010001";
--		WAIT FOR 100 ns;
--				
--		Op <= "0000";--Add_4
--		A <= "10000000000000001100000010100111";
--		B <= "00000000000000000001000000000100";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_5
--		A <= "10000000000000001100000010100111";
--		B <= "10000000000010000001000000000100";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_6
--		-- 15 + 3 = 18
--		A <= "00000000000000000000000000001111";
--		B <= "00000000000000000000000000000011";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_7
--		-- max.no + max.no
--		A <= "01111111111111111111111111111111";
--		B <= "01111111111111111111111111111111";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_8
--		-- max.no + (max.no - 1)
--		A <= "01111111111111111111111111111111";
--		B <= "01111111111111111111111111111110";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_9
--		-- max.no + 1
--		A <= "01111111111111111111111111111111";
--		B <= "00000000000000000000000000000001";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_10
--		-- min.no + min.no
--		A <= "10000000000000000000000000000000";
--		B <= "10000000000000000000000000000000";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_11
--		-- (-1) + (-1)
--		A <= "11111111111111111111111111111111";
--		B <= "11111111111111111111111111111111";
--		WAIT FOR 100 ns;
--		
--		Op <= "0000";--Add_12
--		-- min.no + max.no
--		A <= "11111111111111111111111111111111";
--		B <= "01111111111111111111111111111111";
--		WAIT FOR 100 ns;
		
--		Op <= "0001";--Sub_1
--		-- 0 - 0
--		A <= "00000000000000000000000000000000";
--		B <= "00000000000000000000000000000000";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_2
--		A <= "00000000000000001100000010100111";
--		B <= "00000000000000000001000000000100";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_3
--		A <= "10000000000000001100000010100111";
--		B <= "10000000000010000001000000000100";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_4
--		A <= "00000000000000000000000010100111";
--		B <= "10000000000000000000000000000100";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_4
--		A <= "10000000000000000000000000000100";
--		B <= "00000000000000000000000010100111";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_5
--		-- min.no - min.no
--		A <= "10000000000000000000000000000000";
--		B <= "10000000000000000000000000000000";
--		WAIT FOR 100 ns;
--		
--		-------------- Subtraction -------------
--		Op <= "0001";--Sub_6
--		-- (-1) - (-1)
--		A <= "11111111111111111111111111111111";
--		B <= "11111111111111111111111111111111";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_7
--		-- min.no - max.no
--		A <= "11111111111111111111111111111111";
--		B <= "01111111111111111111111111111111";
--		WAIT FOR 100 ns;
--		
--		Op <= "0001";--Sub_8
--		-- max.no - min.no
--		A <= "01111111111111111111111111111111";
--		B <= "11111111111111111111111111111111";
--		WAIT FOR 100 ns;
		
		------------- AND, OR, NOT -------------
		--------------- NOR, NAND --------------
		Op <= "0010";--AND
		A <= "00000000000000000000000000000111";
		B <= "00000000000000000000000000000100";
		WAIT FOR 100 ns;
		
		Op <= "0010";--AND
		A <= "00100000100001111100010000000111";
		B <= "00100010100001011100010011010100";
		WAIT FOR 100 ns;
		
		Op <= "0011";--OR
		A <= "00000000000000000000000000000111";
		B <= "00000000000000000000000000000100";
		WAIT FOR 100 ns;
		
		Op <= "0011";--OR
		A <= "00100000100001111100010000000111";
		B <= "00100010100001011100010011010100";
		WAIT FOR 100 ns;
		
		Op <= "0100";--NOT
		A <= "00100000100001111100010000000111";
		WAIT FOR 100 ns;
		
		Op <= "0100";--NOT
		A <= "00000000000000000000000000000000";
		WAIT FOR 100 ns;
		
		Op <= "0100";--NOT
		A <= "11111111111111111111111111111111";
		WAIT FOR 100 ns;
		
		Op <= "0110";--NOR
		A <= "00000000000000000000000000000111";
		B <= "00000000000000000000000000000100";
		WAIT FOR 100 ns;
		
		Op <= "0110";--NOR
		A <= "00100000100001111100010000000111";
		B <= "00100010100001011100010011010100";
		WAIT FOR 100 ns;
		
		Op <= "0101";--NAND
		A <= "00000000000000000000000000000111";
		B <= "00000000000000000000000000000100";
		WAIT FOR 100 ns;
		
		Op <= "0101";--NAND
		A <= "00100000100001111100010000000111";
		B <= "00100010100001011100010011010100";
		WAIT FOR 100 ns;
		
		---------------- Shift ----------------
		Op <= "1000";--shift right arithmetic
		A <= "11100000011000000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1000";--shift right arithmetic
		A <= "01111011111110000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1001";--shift right logical
		A <= "11111100000000000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1001";--shift right logical
		A <= "00011110011110000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1010";--shift left logical
		A <= "10000000000000000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1010";--shift left logical
		A <= "10000011111110000000001100001100";
		WAIT FOR 100 ns;
		
		--------------- Rotate ----------------
		Op <= "1100";--rotate left 1
		A <= "10000000000010001000001100000110";
		WAIT FOR 100 ns;
		
		Op <= "1100";--rotate left 1
		A <= "00100011111110000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1101";--rotate right 1
		A <= "00000000000000000000001100000111";
		WAIT FOR 100 ns;
		
		Op <= "1101";--rotate right 1
		A <= "10000011111110000000001100000111";
		WAIT FOR 100 ns;
		WAIT;
	END PROCESS;
END;
-------------------------------------------------------------------------------